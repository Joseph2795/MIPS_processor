`timescale 1ns / 1ps

module mem_inst(
    input wire [4:0] dir,
    input wire [4:0] dir2,
    output reg [31:0] ins,
    output reg [31:0] ins2
    );
    always@*
    begin
        case(dir)
            default:
                ins=32'h00000000;
            5'h00:
                ins=32'h00221803;
            5'h01:
                ins=32'h0C850001;
            5'h02:
                ins=32'h01063804;
            5'h03:
                ins=32'h016C2005;
            5'h04:
                ins=32'h1C090001;
            5'h05:
                ins=32'h0294A007; 
            5'h06:
                ins=32'h01AE7801;
            5'h07:
                ins=32'h06100000;
            5'h08:
                ins=32'h02208806;
            5'h09:
                ins=32'h02529002;
            5'h0A:
                ins=32'h0A730000;
            5'h0B:
                ins=32'h180A0001;
            5'h0C:
                ins=32'h14210001;
            5'h0D:
                ins=32'h00000000;
            5'h0E:
                ins=32'h00000000;
            5'h0F:
                ins=32'h20000014;
            5'h10:
                ins=32'h00000000;
            5'h11:
                ins=32'h00000000;
            5'h12:
                ins=32'h00000000;  
            5'h13:
                ins=32'h00000000;
            5'h14:
                ins=32'h10210000;
            5'h15:
                ins=32'h00000000;
            5'h16:
                ins=32'h00000000;
            5'h17:
                ins=32'h00000000;      
        endcase           
    end  
    always@*
    begin
        case(dir2)
            default:
                ins2=32'h00000000;
            5'h00:
                ins2=32'h00221803;
            5'h01:
                ins2=32'h0C850001;
            5'h02:
                ins2=32'h01063804;
            5'h03:
                ins2=32'h016C2005;
            5'h04:
                ins2=32'h1C090001;
            5'h05:
                ins2=32'h0294A007; 
            5'h06:
                ins2=32'h01AE7801;
            5'h07:
                ins2=32'h06100000;
            5'h08:
                ins2=32'h02208806;
            5'h09:
                ins2=32'h02529002;
            5'h0A:
                ins2=32'h0A730000;
            5'h0B:
                ins2=32'h180A0001;
            5'h0C:
                ins2=32'h14210001;
            5'h0D:
                ins2=32'h00000000;
            5'h0E:
                ins2=32'h00000000;
            5'h0F:
                ins2=32'h20000014;
            5'h10:
                ins2=32'h00000000;
            5'h11:
                ins2=32'h00000000;
            5'h12:
                ins2=32'h00000000;  
            5'h13:
                ins2=32'h00000000;
            5'h14:
                ins2=32'h10210000;
            5'h15:
                ins2=32'h00000000;
            5'h16:
                ins2=32'h00000000;
            5'h17:
                ins2=32'h00000000;
        endcase 
    end
    
endmodule